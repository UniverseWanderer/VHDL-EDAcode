LIBRARY IEEE;--division
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
ENTITY MA IS
PORT(CLK: IN  STD_LOGIC;
	DATA: IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
	FOUT: OUT STD_LOGIC);
END MA;

ARCHITECTURE BEH OF MA IS
	SIGNAL CO,FOUT1,FOUT2	:	STD_LOGIC;
	SIGNAL C1,C2,CLK1,CLK2	:	STD_LOGIC;
	SIGNAL Q1,Q2			: 	STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
	PROCESS(CLK)
	BEGIN
		
		IF (CONV_INTEGER(DATA) REM 2)=1 THEN C1<=CLK;FOUT<=FOUT1;
		ELSIF (CONV_INTEGER(DATA) REM 2)=0 THEN C2<=CLK;FOUT<=FOUT2;
		END IF;
	END PROCESS;
	
	PROCESS(C2)--EVEN
		VARIABLE Q	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	BEGIN
		IF C2'EVENT AND C2='1' THEN
			IF Q<CONV_INTEGER(DATA)/2-1 THEN 
				Q:=Q+1;
			ELSE 
				CO<=NOT(CO);
				Q:=(OTHERS=>'0');
			END IF;
		END IF;
		FOUT2<=CO;
	END PROCESS;
	
	
	PROCESS(C1)--ODD 
	BEGIN
		IF C1'EVENT AND C1='1' THEN 
		  IF(Q1<CONV_INTEGER(DATA)-1) THEN	
			Q1<=Q1+1;
		  ELSE
		    Q1<=(OTHERS=>'0');
		  END IF;
		  IF(Q1<(CONV_INTEGER(DATA)-1)/2) THEN
			CLK1<='1';
		  ELSE 
			CLK1<='0';
		  END IF;
		END IF;
	END PROCESS;
	
	PROCESS(C1)--ODD
	BEGIN
		IF C1'EVENT AND C1='0' THEN
		  IF(Q2<CONV_INTEGER(DATA)-1) THEN	
			Q2<=Q2+1;
		  ELSE
		    Q2<=(OTHERS=>'0');
		  END IF;
		  IF(Q2<(CONV_INTEGER(DATA)-1)/2) THEN
			CLK2<='1';
		  ELSE 
			CLK2<='0';
		  END IF;
		END IF;
	END PROCESS;
	FOUT1<=CLK1 OR CLK2;
	
END BEH;