LIBRARY IEEE;--ODD DIVISION
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY MA IS
PORT(CLK: IN  STD_LOGIC;
	DATA: IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
	FOUT: OUT STD_LOGIC);
END MA;

ARCHITECTURE BEH OF MA IS
	SIGNAL CLK1,CLK2	:	STD_LOGIC;
	SIGNAL Q1,Q2: 	STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
	PROCESS(CLK) 
	BEGIN
		IF CLK'EVENT AND CLK='1' THEN 
		  IF(Q1<CONV_INTEGER(DATA)-1) THEN	
			Q1<=Q1+1;
		  ELSE
		    Q1<=(OTHERS=>'0');
		  END IF;
		  IF(Q1<(CONV_INTEGER(DATA)-1)/2) THEN
			CLK1<='1';
		  ELSE 
			CLK1<='0';
		  END IF;
		END IF;
	END PROCESS;
	
	PROCESS(CLK)
	BEGIN
		IF CLK'EVENT AND CLK='0' THEN
		  IF(Q2<CONV_INTEGER(DATA)-1) THEN	
			Q2<=Q2+1;
		  ELSE
		    Q2<=(OTHERS=>'0');
		  END IF;
		  IF(Q2<(CONV_INTEGER(DATA)-1)/2) THEN
			CLK2<='1';
		  ELSE 
			CLK2<='0';
		  END IF;
		END IF;
	END PROCESS;
	FOUT<=CLK1 OR CLK2;	
END BEH;
