LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY led2 IS
  PORT(CLK,RST,EN   : IN  STD_LOGIC;
	   DEL   		: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
	   LEDAG 		: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END;
ARCHITECTURE bhv OF led2 IS
  BEGIN
	PROCESS(CLK,RST,EN) 
		VARIABLE Q1  : STD_LOGIC_VECTOR(3 DOWNTO 0);
		VARIABLE SEL : STD_LOGIC_VECTOR(2 DOWNTO 0);
		VARIABLE TEMP: INTEGER;
	BEGIN
		IF RST='0' THEN Q1:=(OTHERS=>'0');
		  ELSIF CLK'EVENT AND CLK='1' THEN
			IF TEMP>500 THEN
			  IF EN='1' THEN --start counting
				IF Q1<9 THEN Q1:=Q1+1;
					ELSE Q1:=(OTHERS=>'0');
				END IF;
			  END IF;
			  TEMP:=0;
			ELSE
			  TEMP:=TEMP+1;
			END IF;			
		END IF;

		CASE(Q1) IS
			WHEN "0000" => LEDAG<="0111111";
			WHEN "0001" => LEDAG<="0000110";
			WHEN "0010" => LEDAG<="1011011";
			WHEN "0011" => LEDAG<="1001111";
			WHEN "0100" => LEDAG<="1100110";
			WHEN "0101" => LEDAG<="1101101";
			WHEN "0110" => LEDAG<="1111101";
			WHEN "0111" => LEDAG<="0000111";
			WHEN "1000" => LEDAG<="1111111";
			WHEN "1001" => LEDAG<="1101111";
			WHEN OTHERS => NULL;
		END CASE;
		
		IF CLK'EVENT AND CLK='1' THEN
		    SEL:=SEL+1;		  
		END IF;
		DEL <= SEL;

	END PROCESS;
END bhv;
