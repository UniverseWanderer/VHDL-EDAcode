LIBRARY IEEE;--even division
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY MA IS
PORT(CLK: IN  STD_LOGIC;
	DATA: IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
	FOUT: OUT STD_LOGIC);
END MA;

ARCHITECTURE BEH OF MA IS
	SIGNAL CO	:	STD_LOGIC;
BEGIN
	PROCESS(CLK)
		VARIABLE Q	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	BEGIN
		IF CLK'EVENT AND CLK='1' THEN
			IF Q<CONV_INTEGER(DATA)/2-1 THEN 
				Q:=Q+1;
			ELSE 
				CO<=NOT(CO);
				Q:=(OTHERS=>'0');
			END IF;
		END IF;
		FOUT<=CO;
	END PROCESS;
END BEH;