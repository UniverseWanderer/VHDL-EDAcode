LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY MA IS
PORT(CLK : IN  STD_LOGIC;
	OPT	 : IN  STD_LOGIC;
	RN,CN: OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END MA;

ARCHITECTURE BEH OF MA IS
BEGIN 
	PROCESS(CLK)
		VARIABLE T	: INTEGER RANGE 0 TO 15;
		VARIABLE QR,QC	: STD_LOGIC_VECTOR(15 DOWNTO 0);
	BEGIN
		IF CLK'EVENT AND CLK='1' THEN
		  IF OPT='1' THEN
			IF T<16 THEN				
				CASE(T)IS
					WHEN 0  => QC:="1111111111111110";QR:="0001000000000000";
					WHEN 1  => QC:="1111111111111101";QR:="0111111111111100";
					WHEN 2  => QC:="1111111111111011";QR:="0000000100000000";
					WHEN 3  => QC:="1111111111110111";QR:="0000000100000000";
					WHEN 4  => QC:="1111111111101111";QR:="0000000100000000";
					WHEN 5  => QC:="1111111111011111";QR:="0000000100000000";
					WHEN 6  => QC:="1111111110111111";QR:="0001000100000000";
					WHEN 7  => QC:="1111111101111111";QR:="0011111111111000";
					WHEN 8  => QC:="1111111011111111";QR:="0000000100000000";
					WHEN 9  => QC:="1111110111111111";QR:="0000000100000000";
					WHEN 10 => QC:="1111101111111111";QR:="0000000100000000";
					WHEN 11 => QC:="1111011111111111";QR:="0000000100000000";
					WHEN 12 => QC:="1110111111111111";QR:="0000000100000000";
					WHEN 13 => QC:="1101111111111111";QR:="0010000100000000";
					WHEN 14 => QC:="1011111111111111";QR:="0111111111111111";
					WHEN 15 => QC:="0111111111111111";QR:="0000000000000000";
					WHEN OTHERS => NULL;
				END CASE;				
				T:=T+1;
			ELSE
				T:=0;
			END IF;
		  END IF;
		
		  IF OPT='0' THEN
			IF T<16 THEN				
				CASE(T)IS
					WHEN 0  => QC:="1111111111111110";QR:="0000000001000000";
					WHEN 1  => QC:="1111111111111101";QR:="0000000001000000";
					WHEN 2  => QC:="1111111111111011";QR:="0010000001000000";
					WHEN 3  => QC:="1111111111110111";QR:="0111111111111111";
					WHEN 4  => QC:="1111111111101111";QR:="0000000000100000";
					WHEN 5  => QC:="1111111111011111";QR:="0000000010010000";
					WHEN 6  => QC:="1111111110111111";QR:="0000000010010000";
					WHEN 7  => QC:="1111111101111111";QR:="0000100010001000";
					WHEN 8  => QC:="1111111011111111";QR:="0001111111111100";
					WHEN 9  => QC:="1111110111111111";QR:="0000000010000000";
					WHEN 10 => QC:="1111101111111111";QR:="0000001010010000";
					WHEN 11 => QC:="1111011111111111";QR:="0000010010010000";
					WHEN 12 => QC:="1110111111111111";QR:="0000100010001000";
					WHEN 13 => QC:="1101111111111111";QR:="0001100010000100";
					WHEN 14 => QC:="1011111111111111";QR:="0001000010100010";
					WHEN 15 => QC:="0111111111111111";QR:="0000000001000000";
					WHEN OTHERS => NULL;
				END CASE;				
				T:=T+1;
			ELSE
				T:=0;
			END IF;
		  END IF;
												
		END IF;
		CN<=QR; 
		RN<=QC;		
	END PROCESS;
END BEH;