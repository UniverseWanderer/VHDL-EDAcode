LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY exp2 IS
  PORT(K : IN  STD_LOGIC_VECTOR(11 DOWNTO 0);
	   D : OUT STD_LOGIC_VECTOR(11 DOWNTO 0));
END;

ARCHITECTURE bhv OF exp2 IS
  BEGIN
	PROCESS(K) BEGIN
	D(11)<=K(11);
DO: FOR n IN 1 TO 11 LOOP
	D(11-n)<=K(11-n) XOR K(12-n);
	END LOOP DO;
	END PROCESS;
END;